
module altpll (
	clk_clk,
	clock_30_clk,
	reset_reset_n);	

	input		clk_clk;
	output		clock_30_clk;
	input		reset_reset_n;
endmodule
