module NumberDecoder(
    input clk, 
    input rst_n,

    input [17:0] i_data,
    output [31:0] o_seven
);

logic [31:0] n_o_seven;

logic [17:0] temp [0:6];
endmodule