`ifdef PEARRAY
`else
`define PEARRAY

`include "util.v"

module PEArray (
	input clk,    // Clock
	input rst_n,  // Asynchronous reset active low
	
);

endmodule
`endif